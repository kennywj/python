//The Netlist from Uncle 
module ncl_mac ( rst_n  ,  t_ina  ,  f_ina  ,  t_inb  ,  f_inb  ,  t_coef  ,  f_coef  ,  t_mac_out  ,  f_mac_out  , 
 ackout  ,  ackin );
  input ackin ;
  output ackout ;
  output [7:0] f_mac_out ;
  output [7:0] t_mac_out ;
  input [3:0] f_coef ;
  input [3:0] t_coef ;
  input [3:0] f_inb ;
  input [3:0] t_inb ;
  input [3:0] f_ina ;
  input [3:0] t_ina ;
  input rst_n ;
  wire [3:0] f_ina_reg ;
  wire [3:0] t_ina_reg ;
  wire [3:0] f_inb_reg ;
  wire [3:0] t_inb_reg ;
  wire [3:0] f_coef_reg ;
  wire [3:0] t_coef_reg ;
  wire [4:0] f_shift2_reg ;
  wire [4:0] t_shift2_reg ;
  wire [7:0] f_mul_reg ;
  wire [7:0] t_mul_reg ;
  wire acknet42 ;
  wire acknet41 ;
  wire acknet40 ;
  wire acknet39 ;
  wire acknet38 ;
  wire acknet37 ;
  wire acknet36 ;
  wire acknet35 ;
  wire acknet34 ;
  wire acknet33 ;
  wire acknet32 ;
  wire acknet31 ;
  wire acknet30 ;
  wire acknet29 ;
  wire acknet28 ;
  wire acknet27 ;
  wire acknet26 ;
  wire acknet25 ;
  wire acknet24 ;
  wire acknet23 ;
  wire acknet22 ;
  wire acknet21 ;
  wire acknet20 ;
  wire acknet19 ;
  wire acknet18 ;
  wire acknet17 ;
  wire acknet16 ;
  wire acknet15 ;
  wire acknet14 ;
  wire acknet13 ;
  wire acknet12 ;
  wire acknet11 ;
  wire acknet10 ;
  wire acknet9 ;
  wire acknet8 ;
  wire acknet7 ;
  wire acknet6 ;
  wire acknet5 ;
  wire acknet4 ;
  wire acknet3 ;
  wire acknet2 ;
  wire acknet1 ;
  wire acknet0 ;
  wire f_n37 ;
  wire t_n37 ;
  wire f_n36 ;
  wire t_n36 ;
  wire f_n40 ;
  wire t_n40 ;
  wire f_n39 ;
  wire t_n39 ;
  wire f_n38 ;
  wire t_n38 ;
  wire f_n41 ;
  wire t_n41 ;
  wire f_n43 ;
  wire t_n43 ;
  wire f_n42 ;
  wire t_n42 ;
  wire f_n45 ;
  wire t_n45 ;
  wire f_n44 ;
  wire t_n44 ;
  wire f_n48 ;
  wire t_n48 ;
  wire f_n47 ;
  wire t_n47 ;
  wire f_n46 ;
  wire t_n46 ;
  wire f_n50 ;
  wire t_n50 ;
  wire f_n49 ;
  wire t_n49 ;
  wire f_n52 ;
  wire t_n52 ;
  wire f_n51 ;
  wire t_n51 ;
  wire f_n53 ;
  wire t_n53 ;
  wire f_N8 ;
  wire t_N8 ;
  wire f_n56 ;
  wire t_n56 ;
  wire f_n54 ;
  wire t_n54 ;
  wire f_N7 ;
  wire t_N7 ;
  wire f_n59 ;
  wire t_n59 ;
  wire f_n58 ;
  wire t_n58 ;
  wire f_n55 ;
  wire t_n55 ;
  wire f_N6 ;
  wire t_N6 ;
  wire f_n62 ;
  wire t_n62 ;
  wire f_n61 ;
  wire t_n61 ;
  wire f_n57 ;
  wire t_n57 ;
  wire f_N5 ;
  wire t_N5 ;
  wire f_n65 ;
  wire t_n65 ;
  wire f_n63 ;
  wire t_n63 ;
  wire f_n60 ;
  wire t_n60 ;
  wire f_N4 ;
  wire t_N4 ;
  wire f_n68 ;
  wire t_n68 ;
  wire f_n67 ;
  wire t_n67 ;
  wire f_n66 ;
  wire t_n66 ;
  wire f_n64 ;
  wire t_n64 ;
  wire f_N3 ;
  wire t_N3 ;
  wire f_N1 ;
  wire t_N1 ;
  wire f_n70 ;
  wire t_n70 ;
  wire f_n69 ;
  wire t_n69 ;
  wire f_N2 ;
  wire t_N2 ;
  wire f_N12 ;
  wire t_N12 ;
  wire f_n71 ;
  wire t_n71 ;
  wire f_N11 ;
  wire t_N11 ;
  wire f_n73 ;
  wire t_n73 ;
  wire f_n72 ;
  wire t_n72 ;
  wire f_N10 ;
  wire t_N10 ;
  wire f_N9 ;
  wire t_N9 ;
  wire f_n74 ;
  wire t_n74 ;
  wire f_N13 ;
  wire t_N13 ;
  wire f_n75 ;
  wire t_n75 ;
  wire f_N14 ;
  wire t_N14 ;
  wire f_n76 ;
  wire t_n76 ;
  wire f_N15 ;
  wire t_N15 ;
  wire f_n77 ;
  wire t_n77 ;
  wire f_N16 ;
  wire t_N16 ;
  wire f_constnet0 ;
  wire t_constnet0 ;
  wire f_n1_N ;
  wire t_n1_N ;
  wire f_n1_N_0 ;
  wire t_n1_N_0 ;
  wire f_n1_N_1 ;
  wire t_n1_N_1 ;
  wire f_n1_N_2 ;
  wire t_n1_N_2 ;
  wire f_q2_N ;
  wire t_q2_N ;
  wire n2_N ;
  wire f_q1_N ;
  wire t_q1_N ;
  wire n1_N ;
  wire f_q2_N_0 ;
  wire t_q2_N_0 ;
  wire n2_N_0 ;
  wire f_q1_N_0 ;
  wire t_q1_N_0 ;
  wire n1_N_0 ;
  wire f_q2_N_1 ;
  wire t_q2_N_1 ;
  wire n2_N_1 ;
  wire f_q1_N_1 ;
  wire t_q1_N_1 ;
  wire n1_N_1 ;
  wire f_q2_N_2 ;
  wire t_q2_N_2 ;
  wire n2_N_2 ;
  wire f_q1_N_2 ;
  wire t_q1_N_2 ;
  wire n1_N_2 ;
  wire f_q2_N_3 ;
  wire t_q2_N_3 ;
  wire n2_N_3 ;
  wire f_q1_N_3 ;
  wire t_q1_N_3 ;
  wire n1_N_3 ;
  wire f_q2_N_4 ;
  wire t_q2_N_4 ;
  wire n2_N_4 ;
  wire f_q1_N_4 ;
  wire t_q1_N_4 ;
  wire n1_N_4 ;
  wire f_q2_N_5 ;
  wire t_q2_N_5 ;
  wire n2_N_5 ;
  wire f_q1_N_5 ;
  wire t_q1_N_5 ;
  wire n1_N_5 ;
  wire f_q2_N_6 ;
  wire t_q2_N_6 ;
  wire n2_N_6 ;
  wire f_q1_N_6 ;
  wire t_q1_N_6 ;
  wire n1_N_6 ;
  wire f_q2_N_7 ;
  wire t_q2_N_7 ;
  wire n2_N_7 ;
  wire f_q1_N_7 ;
  wire t_q1_N_7 ;
  wire n1_N_7 ;
  wire f_q2_N_8 ;
  wire t_q2_N_8 ;
  wire n2_N_8 ;
  wire f_q1_N_8 ;
  wire t_q1_N_8 ;
  wire n1_N_8 ;
  wire f_q2_N_9 ;
  wire t_q2_N_9 ;
  wire n2_N_9 ;
  wire f_q1_N_9 ;
  wire t_q1_N_9 ;
  wire n1_N_9 ;
  wire f_q2_N_10 ;
  wire t_q2_N_10 ;
  wire n2_N_10 ;
  wire f_q1_N_10 ;
  wire t_q1_N_10 ;
  wire n1_N_10 ;
  wire f_q2_N_11 ;
  wire t_q2_N_11 ;
  wire n2_N_11 ;
  wire f_q1_N_11 ;
  wire t_q1_N_11 ;
  wire n1_N_11 ;
  wire f_q2_N_12 ;
  wire t_q2_N_12 ;
  wire n2_N_12 ;
  wire f_q1_N_12 ;
  wire t_q1_N_12 ;
  wire n1_N_12 ;
  wire f_q2_N_13 ;
  wire t_q2_N_13 ;
  wire n2_N_13 ;
  wire f_q1_N_13 ;
  wire t_q1_N_13 ;
  wire n1_N_13 ;
  wire f_q2_N_14 ;
  wire t_q2_N_14 ;
  wire n2_N_14 ;
  wire f_q1_N_14 ;
  wire t_q1_N_14 ;
  wire n1_N_14 ;
  wire f_q2_N_15 ;
  wire t_q2_N_15 ;
  wire n2_N_15 ;
  wire f_q1_N_15 ;
  wire t_q1_N_15 ;
  wire n1_N_15 ;
  wire f_q2_N_16 ;
  wire t_q2_N_16 ;
  wire n2_N_16 ;
  wire f_q1_N_16 ;
  wire t_q1_N_16 ;
  wire n1_N_16 ;
  wire f_q2_N_17 ;
  wire t_q2_N_17 ;
  wire n2_N_17 ;
  wire f_q1_N_17 ;
  wire t_q1_N_17 ;
  wire n1_N_17 ;
  wire f_q2_N_18 ;
  wire t_q2_N_18 ;
  wire n2_N_18 ;
  wire f_q1_N_18 ;
  wire t_q1_N_18 ;
  wire n1_N_18 ;
  wire f_q2_N_19 ;
  wire t_q2_N_19 ;
  wire n2_N_19 ;
  wire f_q1_N_19 ;
  wire t_q1_N_19 ;
  wire n1_N_19 ;
  wire f_q2_N_20 ;
  wire t_q2_N_20 ;
  wire n2_N_20 ;
  wire f_q1_N_20 ;
  wire t_q1_N_20 ;
  wire n1_N_20 ;
  wire f_q2_N_21 ;
  wire t_q2_N_21 ;
  wire n2_N_21 ;
  wire f_q1_N_21 ;
  wire t_q1_N_21 ;
  wire n1_N_21 ;
  wire f_q2_N_22 ;
  wire t_q2_N_22 ;
  wire n2_N_22 ;
  wire f_q1_N_22 ;
  wire t_q1_N_22 ;
  wire n1_N_22 ;
  wire f_q2_N_23 ;
  wire t_q2_N_23 ;
  wire n2_N_23 ;
  wire f_q1_N_23 ;
  wire t_q1_N_23 ;
  wire n1_N_23 ;
  wire f_q2_N_24 ;
  wire t_q2_N_24 ;
  wire n2_N_24 ;
  wire f_q1_N_24 ;
  wire t_q1_N_24 ;
  wire n1_N_24 ;
  wire f_q2_N_25 ;
  wire t_q2_N_25 ;
  wire n2_N_25 ;
  wire f_q1_N_25 ;
  wire t_q1_N_25 ;
  wire n1_N_25 ;
  wire f_q2_N_26 ;
  wire t_q2_N_26 ;
  wire n2_N_26 ;
  wire f_q1_N_26 ;
  wire t_q1_N_26 ;
  wire n1_N_26 ;
  wire f_q2_N_27 ;
  wire t_q2_N_27 ;
  wire n2_N_27 ;
  wire f_q1_N_27 ;
  wire t_q1_N_27 ;
  wire n1_N_27 ;
  wire f_q2_N_28 ;
  wire t_q2_N_28 ;
  wire n2_N_28 ;
  wire f_q1_N_28 ;
  wire t_q1_N_28 ;
  wire n1_N_28 ;
  wire f_q2_N_29 ;
  wire t_q2_N_29 ;
  wire n2_N_29 ;
  wire f_q1_N_29 ;
  wire t_q1_N_29 ;
  wire n1_N_29 ;
  wire f_q2_N_30 ;
  wire t_q2_N_30 ;
  wire n2_N_30 ;
  wire f_q1_N_30 ;
  wire t_q1_N_30 ;
  wire n1_N_30 ;
  wire f_q2_N_31 ;
  wire t_q2_N_31 ;
  wire n2_N_31 ;
  wire f_q1_N_31 ;
  wire t_q1_N_31 ;
  wire n1_N_31 ;
  wire bufnet ;
  wire bufnet_0 ;
  wire bufnet_1 ;
  wire bufnet_2 ;
  wire rst_n ;
  wire ackout ;
  wire ackin ;
  assign ackout = acknet42 ; 
  th23  U52_U_U_2 (.a ( f_n38 ) , .b ( f_n40 ) , .c ( f_n39 ) , .y ( f_n58 ));
  th23  U52_U_U_1 (.a ( t_n38 ) , .b ( t_n40 ) , .c ( t_n39 ) , .y ( t_n58 ));
  th34w2  U52_U_U_0 (.a ( t_n58 ) , .b ( f_n38 ) , .c ( f_n40 ) , .d ( f_n39 ) , .y ( f_n62 ));
  th34w2  U52_U_U (.a ( f_n58 ) , .b ( t_n38 ) , .c ( t_n40 ) , .d ( t_n39 ) , .y ( t_n62 ));
  th23  U72_U_U_2 (.a ( f_n57 ) , .b ( f_n59 ) , .c ( f_n58 ) , .y ( f_n55 ));
  th23  U72_U_U_1 (.a ( t_n57 ) , .b ( t_n59 ) , .c ( t_n58 ) , .y ( t_n55 ));
  th34w2  U72_U_U_0 (.a ( t_n55 ) , .b ( f_n57 ) , .c ( f_n59 ) , .d ( f_n58 ) , .y ( f_N6 ));
  th34w2  U72_U_U (.a ( f_n55 ) , .b ( t_n57 ) , .c ( t_n59 ) , .d ( t_n58 ) , .y ( t_N6 ));
  th23  U73_U_U_2 (.a ( f_n60 ) , .b ( f_n62 ) , .c ( f_n61 ) , .y ( f_n57 ));
  th23  U73_U_U_1 (.a ( t_n60 ) , .b ( t_n62 ) , .c ( t_n61 ) , .y ( t_n57 ));
  th34w2  U73_U_U_0 (.a ( t_n57 ) , .b ( f_n60 ) , .c ( f_n62 ) , .d ( f_n61 ) , .y ( f_N5 ));
  th34w2  U73_U_U (.a ( f_n57 ) , .b ( t_n60 ) , .c ( t_n62 ) , .d ( t_n61 ) , .y ( t_N5 ));
  th23  U74_U_U_2 (.a ( f_n63 ) , .b ( f_n65 ) , .c ( f_n64 ) , .y ( f_n60 ));
  th23  U74_U_U_1 (.a ( t_n63 ) , .b ( t_n65 ) , .c ( t_n64 ) , .y ( t_n60 ));
  th34w2  U74_U_U_0 (.a ( t_n60 ) , .b ( f_n63 ) , .c ( f_n65 ) , .d ( f_n64 ) , .y ( f_N4 ));
  th34w2  U74_U_U (.a ( f_n60 ) , .b ( t_n63 ) , .c ( t_n65 ) , .d ( t_n64 ) , .y ( t_N4 ));
  th23  U75_U_U_2 (.a ( f_n66 ) , .b ( f_n68 ) , .c ( f_n67 ) , .y ( f_n64 ));
  th23  U75_U_U_1 (.a ( t_n66 ) , .b ( t_n68 ) , .c ( t_n67 ) , .y ( t_n64 ));
  th34w2  U75_U_U_0 (.a ( t_n64 ) , .b ( f_n66 ) , .c ( f_n68 ) , .d ( f_n67 ) , .y ( f_N3 ));
  th34w2  U75_U_U (.a ( f_n64 ) , .b ( t_n66 ) , .c ( t_n68 ) , .d ( t_n67 ) , .y ( t_N3 ));
  th23  U79_U_U_2 (.a ( f_n71 ) , .b ( f_mul_reg[3] ) , .c ( f_shift2_reg[3] ) , .y ( f_n74 ));
  th23  U79_U_U_1 (.a ( t_n71 ) , .b ( t_mul_reg[3] ) , .c ( t_shift2_reg[3] ) , .y ( t_n74 ));
  th34w2  U79_U_U_0 (.a ( t_n74 ) , .b ( f_n71 ) , .c ( f_mul_reg[3] ) , .d ( f_shift2_reg[3] ) , .y ( f_N12 ));
  th34w2  U79_U_U (.a ( f_n74 ) , .b ( t_n71 ) , .c ( t_mul_reg[3] ) , .d ( t_shift2_reg[3] ) , .y ( t_N12 ));
  th23  U80_U_U_2 (.a ( f_n72 ) , .b ( f_mul_reg[2] ) , .c ( f_shift2_reg[2] ) , .y ( f_n71 ));
  th23  U80_U_U_1 (.a ( t_n72 ) , .b ( t_mul_reg[2] ) , .c ( t_shift2_reg[2] ) , .y ( t_n71 ));
  th34w2  U80_U_U_0 (.a ( t_n71 ) , .b ( f_n72 ) , .c ( f_mul_reg[2] ) , .d ( f_shift2_reg[2] ) , .y ( f_N11 ));
  th34w2  U80_U_U (.a ( f_n71 ) , .b ( t_n72 ) , .c ( t_mul_reg[2] ) , .d ( t_shift2_reg[2] ) , .y ( t_N11 ));
  th23  U81_U_U_2 (.a ( f_n73 ) , .b ( f_mul_reg[1] ) , .c ( f_shift2_reg[1] ) , .y ( f_n72 ));
  th23  U81_U_U_1 (.a ( t_n73 ) , .b ( t_mul_reg[1] ) , .c ( t_shift2_reg[1] ) , .y ( t_n72 ));
  th34w2  U81_U_U_0 (.a ( t_n72 ) , .b ( f_n73 ) , .c ( f_mul_reg[1] ) , .d ( f_shift2_reg[1] ) , .y ( f_N10 ));
  th34w2  U81_U_U (.a ( f_n72 ) , .b ( t_n73 ) , .c ( t_mul_reg[1] ) , .d ( t_shift2_reg[1] ) , .y ( t_N10 ));
  th23  U83_U_U_2 (.a ( f_n74 ) , .b ( f_mul_reg[4] ) , .c ( f_shift2_reg[4] ) , .y ( f_n75 ));
  th23  U83_U_U_1 (.a ( t_n74 ) , .b ( t_mul_reg[4] ) , .c ( t_shift2_reg[4] ) , .y ( t_n75 ));
  th34w2  U83_U_U_0 (.a ( t_n75 ) , .b ( f_n74 ) , .c ( f_mul_reg[4] ) , .d ( f_shift2_reg[4] ) , .y ( f_N13 ));
  th34w2  U83_U_U (.a ( f_n75 ) , .b ( t_n74 ) , .c ( t_mul_reg[4] ) , .d ( t_shift2_reg[4] ) , .y ( t_N13 ));
  th23  U84_U_U_2 (.a ( f_n75 ) , .b ( f_mul_reg[5] ) , .c ( f_shift2_reg[0] ) , .y ( f_n76 ));
  th23  U84_U_U_1 (.a ( t_n75 ) , .b ( t_mul_reg[5] ) , .c ( t_shift2_reg[0] ) , .y ( t_n76 ));
  th34w2  U84_U_U_0 (.a ( t_n76 ) , .b ( f_n75 ) , .c ( f_mul_reg[5] ) , .d ( f_shift2_reg[0] ) , .y ( f_N14 ));
  th34w2  U84_U_U (.a ( f_n76 ) , .b ( t_n75 ) , .c ( t_mul_reg[5] ) , .d ( t_shift2_reg[0] ) , .y ( t_N14 ));
  th23  U85_U_U_2 (.a ( f_n76 ) , .b ( f_mul_reg[6] ) , .c ( f_shift2_reg[0] ) , .y ( f_n77 ));
  th23  U85_U_U_1 (.a ( t_n76 ) , .b ( t_mul_reg[6] ) , .c ( t_shift2_reg[0] ) , .y ( t_n77 ));
  th34w2  U85_U_U_0 (.a ( t_n77 ) , .b ( f_n76 ) , .c ( f_mul_reg[6] ) , .d ( f_shift2_reg[0] ) , .y ( f_N15 ));
  th34w2  U85_U_U (.a ( f_n77 ) , .b ( t_n76 ) , .c ( t_mul_reg[6] ) , .d ( t_shift2_reg[0] ) , .y ( t_N15 ));
  th33  cgate9 (.a ( acknet41 ) , .b ( acknet40 ) , .c ( acknet39 ) , .y ( acknet42 ));
  th44  cgate8 (.a ( acknet26 ) , .b ( acknet29 ) , .c ( acknet32 ) , .d ( acknet21 ) , .y ( acknet41 ));
  th44  cgate7 (.a ( acknet25 ) , .b ( acknet28 ) , .c ( acknet31 ) , .d ( acknet23 ) , .y ( acknet40 ));
  th44  cgate6 (.a ( acknet24 ) , .b ( acknet27 ) , .c ( acknet30 ) , .d ( acknet22 ) , .y ( acknet39 ));
  th22  cgate5 (.a ( acknet37 ) , .b ( acknet36 ) , .y ( acknet38 ));
  th44  cgate4 (.a ( acknet7 ) , .b ( acknet2 ) , .c ( acknet5 ) , .d ( acknet8 ) , .y ( acknet37 ));
  th44  cgate3 (.a ( acknet3 ) , .b ( acknet6 ) , .c ( acknet1 ) , .d ( acknet4 ) , .y ( acknet36 ));
  th22  cgate2 (.a ( acknet34 ) , .b ( acknet33 ) , .y ( acknet35 ));
  th44  cgate1 (.a ( acknet13 ) , .b ( acknet20 ) , .c ( acknet15 ) , .d ( acknet18 ) , .y ( acknet34 ));
  th44  cgate0 (.a ( acknet16 ) , .b ( acknet19 ) , .c ( acknet14 ) , .d ( acknet17 ) , .y ( acknet33 ));
  th24comp  U82_U (.y ( t_N9 ) , .d ( f_shift2_reg[0] ) , .c ( f_mul_reg[0] ) , .b ( t_mul_reg[0] ) , .a ( t_shift2_reg[0] ));
  th24comp  U82_U_0 (.y ( f_N9 ) , .d ( f_shift2_reg[0] ) , .c ( t_mul_reg[0] ) , .b ( f_mul_reg[0] ) , .a ( t_shift2_reg[0] ));
  thand0  U78_U (.y ( f_n73 ) , .d ( t_mul_reg[0] ) , .c ( t_shift2_reg[0] ) , .b ( f_mul_reg[0] ) , .a ( f_shift2_reg[0] ));
  th22  U78_U_0 (.y ( t_n73 ) , .b ( t_mul_reg[0] ) , .a ( t_shift2_reg[0] ));
  th24comp  U77_U (.y ( t_N2 ) , .d ( f_n70 ) , .c ( f_n69 ) , .b ( t_n69 ) , .a ( t_n70 ));
  th24comp  U77_U_0 (.y ( f_N2 ) , .d ( f_n70 ) , .c ( t_n69 ) , .b ( f_n69 ) , .a ( t_n70 ));
  thand0  U76_U (.y ( f_N1 ) , .d ( t_inb_reg[0] ) , .c ( t_ina_reg[0] ) , .b ( f_inb_reg[0] ) , .a ( f_ina_reg[0] ));
  th22  U76_U_0 (.y ( t_N1 ) , .b ( t_inb_reg[0] ) , .a ( t_ina_reg[0] ));
  thand0  U70_U (.y ( f_N8 ) , .d ( t_n53 ) , .c ( t_n56 ) , .b ( f_n53 ) , .a ( f_n56 ));
  th22  U70_U_0 (.y ( t_N8 ) , .b ( t_n53 ) , .a ( t_n56 ));
  thand0  U69_U (.y ( t_n53 ) , .d ( f_n54 ) , .c ( f_n55 ) , .b ( t_n54 ) , .a ( t_n55 ));
  th22  U69_U_0 (.y ( f_n53 ) , .b ( f_n54 ) , .a ( f_n55 ));
  thand0  U68_U (.y ( t_n54 ) , .d ( f_n51 ) , .c ( f_n52 ) , .b ( t_n51 ) , .a ( t_n52 ));
  th22  U68_U_0 (.y ( f_n54 ) , .b ( f_n51 ) , .a ( f_n52 ));
  thand0  U67_U (.y ( f_n51 ) , .d ( t_n49 ) , .c ( t_n50 ) , .b ( f_n49 ) , .a ( f_n50 ));
  th22  U67_U_0 (.y ( t_n51 ) , .b ( t_n49 ) , .a ( t_n50 ));
  thand0  U65_U (.y ( f_n66 ) , .d ( t_inb_reg[0] ) , .c ( t_ina_reg[2] ) , .b ( f_inb_reg[0] ) , .a ( f_ina_reg[2] ));
  th22  U65_U_0 (.y ( t_n66 ) , .b ( t_inb_reg[0] ) , .a ( t_ina_reg[2] ));
  thand0  U64_U (.y ( f_n67 ) , .d ( t_n69 ) , .c ( t_n70 ) , .b ( f_n69 ) , .a ( f_n70 ));
  th22  U64_U_0 (.y ( t_n67 ) , .b ( t_n69 ) , .a ( t_n70 ));
  thand0  U63_U (.y ( f_n69 ) , .d ( t_inb_reg[0] ) , .c ( t_ina_reg[1] ) , .b ( f_inb_reg[0] ) , .a ( f_ina_reg[1] ));
  th22  U63_U_0 (.y ( t_n69 ) , .b ( t_inb_reg[0] ) , .a ( t_ina_reg[1] ));
  thand0  U62_U (.y ( f_n70 ) , .d ( t_ina_reg[0] ) , .c ( t_inb_reg[1] ) , .b ( f_ina_reg[0] ) , .a ( f_inb_reg[1] ));
  th22  U62_U_0 (.y ( t_n70 ) , .b ( t_ina_reg[0] ) , .a ( t_inb_reg[1] ));
  th24comp  U61_U (.y ( t_n68 ) , .d ( f_n45 ) , .c ( f_n44 ) , .b ( t_n44 ) , .a ( t_n45 ));
  th24comp  U61_U_0 (.y ( f_n68 ) , .d ( f_n45 ) , .c ( t_n44 ) , .b ( f_n44 ) , .a ( t_n45 ));
  th24comp  U60_U (.y ( t_n65 ) , .d ( f_n43 ) , .c ( f_n42 ) , .b ( t_n42 ) , .a ( t_n43 ));
  th24comp  U60_U_0 (.y ( f_n65 ) , .d ( f_n43 ) , .c ( t_n42 ) , .b ( f_n42 ) , .a ( t_n43 ));
  thand0  U59_U (.y ( t_n61 ) , .d ( f_n41 ) , .c ( f_n48 ) , .b ( t_n41 ) , .a ( t_n48 ));
  th22  U59_U_0 (.y ( f_n61 ) , .b ( f_n41 ) , .a ( f_n48 ));
  thand0  U58_U (.y ( f_n41 ) , .d ( t_n47 ) , .c ( t_n46 ) , .b ( f_n47 ) , .a ( f_n46 ));
  th22  U58_U_0 (.y ( t_n41 ) , .b ( t_n47 ) , .a ( t_n46 ));
  thand0  U57_U (.y ( f_n47 ) , .d ( t_inb_reg[0] ) , .c ( t_ina_reg[3] ) , .b ( f_inb_reg[0] ) , .a ( f_ina_reg[3] ));
  th22  U57_U_0 (.y ( t_n47 ) , .b ( t_inb_reg[0] ) , .a ( t_ina_reg[3] ));
  thand0  U56_U (.y ( f_n46 ) , .d ( t_ina_reg[1] ) , .c ( t_inb_reg[2] ) , .b ( f_ina_reg[1] ) , .a ( f_inb_reg[2] ));
  th22  U56_U_0 (.y ( t_n46 ) , .b ( t_ina_reg[1] ) , .a ( t_inb_reg[2] ));
  thand0  U55_U (.y ( f_n48 ) , .d ( t_n44 ) , .c ( t_n45 ) , .b ( f_n44 ) , .a ( f_n45 ));
  th22  U55_U_0 (.y ( t_n48 ) , .b ( t_n44 ) , .a ( t_n45 ));
  thand0  U54_U (.y ( f_n44 ) , .d ( t_ina_reg[0] ) , .c ( t_inb_reg[2] ) , .b ( f_ina_reg[0] ) , .a ( f_inb_reg[2] ));
  th22  U54_U_0 (.y ( t_n44 ) , .b ( t_ina_reg[0] ) , .a ( t_inb_reg[2] ));
  thand0  U53_U (.y ( f_n45 ) , .d ( t_inb_reg[1] ) , .c ( t_ina_reg[1] ) , .b ( f_inb_reg[1] ) , .a ( f_ina_reg[1] ));
  th22  U53_U_0 (.y ( t_n45 ) , .b ( t_inb_reg[1] ) , .a ( t_ina_reg[1] ));
  thand0  U51_U (.y ( f_n38 ) , .d ( t_inb_reg[1] ) , .c ( t_ina_reg[3] ) , .b ( f_inb_reg[1] ) , .a ( f_ina_reg[3] ));
  th22  U51_U_0 (.y ( t_n38 ) , .b ( t_inb_reg[1] ) , .a ( t_ina_reg[3] ));
  thand0  U50_U (.y ( f_n39 ) , .d ( t_n42 ) , .c ( t_n43 ) , .b ( f_n42 ) , .a ( f_n43 ));
  th22  U50_U_0 (.y ( t_n39 ) , .b ( t_n42 ) , .a ( t_n43 ));
  thand0  U49_U (.y ( f_n42 ) , .d ( t_inb_reg[1] ) , .c ( t_ina_reg[2] ) , .b ( f_inb_reg[1] ) , .a ( f_ina_reg[2] ));
  th22  U49_U_0 (.y ( t_n42 ) , .b ( t_inb_reg[1] ) , .a ( t_ina_reg[2] ));
  thand0  U48_U (.y ( f_n43 ) , .d ( t_ina_reg[0] ) , .c ( t_inb_reg[3] ) , .b ( f_ina_reg[0] ) , .a ( f_inb_reg[3] ));
  th22  U48_U_0 (.y ( t_n43 ) , .b ( t_ina_reg[0] ) , .a ( t_inb_reg[3] ));
  th24comp  U47_U (.y ( t_n40 ) , .d ( f_n37 ) , .c ( f_n36 ) , .b ( t_n36 ) , .a ( t_n37 ));
  th24comp  U47_U_0 (.y ( f_n40 ) , .d ( f_n37 ) , .c ( t_n36 ) , .b ( f_n36 ) , .a ( t_n37 ));
  thand0  U45_U (.y ( f_n49 ) , .d ( t_ina_reg[2] ) , .c ( t_inb_reg[3] ) , .b ( f_ina_reg[2] ) , .a ( f_inb_reg[3] ));
  th22  U45_U_0 (.y ( t_n49 ) , .b ( t_ina_reg[2] ) , .a ( t_inb_reg[3] ));
  thand0  U44_U (.y ( f_n50 ) , .d ( t_inb_reg[2] ) , .c ( t_ina_reg[3] ) , .b ( f_inb_reg[2] ) , .a ( f_ina_reg[3] ));
  th22  U44_U_0 (.y ( t_n50 ) , .b ( t_inb_reg[2] ) , .a ( t_ina_reg[3] ));
  thand0  U43_U (.y ( f_n52 ) , .d ( t_n36 ) , .c ( t_n37 ) , .b ( f_n36 ) , .a ( f_n37 ));
  th22  U43_U_0 (.y ( t_n52 ) , .b ( t_n36 ) , .a ( t_n37 ));
  thand0  U42_U (.y ( f_n36 ) , .d ( t_ina_reg[1] ) , .c ( t_inb_reg[3] ) , .b ( f_ina_reg[1] ) , .a ( f_inb_reg[3] ));
  th22  U42_U_0 (.y ( t_n36 ) , .b ( t_ina_reg[1] ) , .a ( t_inb_reg[3] ));
  thand0  U41_U (.y ( f_n37 ) , .d ( t_ina_reg[2] ) , .c ( t_inb_reg[2] ) , .b ( f_ina_reg[2] ) , .a ( f_inb_reg[2] ));
  th22  U41_U_0 (.y ( t_n37 ) , .b ( t_ina_reg[2] ) , .a ( t_inb_reg[2] ));
  thand0  U40_U (.y ( f_n56 ) , .d ( t_ina_reg[3] ) , .c ( t_inb_reg[3] ) , .b ( f_ina_reg[3] ) , .a ( f_inb_reg[3] ));
  th22  U40_U_0 (.y ( t_n56 ) , .b ( t_ina_reg[3] ) , .a ( t_inb_reg[3] ));
  th24comp  U46_U_0_U (.y ( t_n1_N_2 ) , .d ( f_n52 ) , .c ( f_n50 ) , .b ( t_n50 ) , .a ( t_n52 ));
  th24comp  U46_U_0_U_0 (.y ( f_n1_N_2 ) , .d ( f_n52 ) , .c ( t_n50 ) , .b ( f_n50 ) , .a ( t_n52 ));
  th24comp  U46_U_U (.y ( t_n59 ) , .d ( f_n1_N_2 ) , .c ( f_n49 ) , .b ( t_n49 ) , .a ( t_n1_N_2 ));
  th24comp  U46_U_U_0 (.y ( f_n59 ) , .d ( f_n1_N_2 ) , .c ( t_n49 ) , .b ( f_n49 ) , .a ( t_n1_N_2 ));
  th24comp  U66_U_0_U (.y ( t_n1_N_1 ) , .d ( f_n48 ) , .c ( f_n47 ) , .b ( t_n47 ) , .a ( t_n48 ));
  th24comp  U66_U_0_U_0 (.y ( f_n1_N_1 ) , .d ( f_n48 ) , .c ( t_n47 ) , .b ( f_n47 ) , .a ( t_n48 ));
  th24comp  U66_U_U (.y ( t_n63 ) , .d ( f_n1_N_1 ) , .c ( f_n46 ) , .b ( t_n46 ) , .a ( t_n1_N_1 ));
  th24comp  U66_U_U_0 (.y ( f_n63 ) , .d ( f_n1_N_1 ) , .c ( t_n46 ) , .b ( f_n46 ) , .a ( t_n1_N_1 ));
  th24comp  U71_U_0_U (.y ( t_n1_N_0 ) , .d ( f_n56 ) , .c ( f_n55 ) , .b ( t_n55 ) , .a ( t_n56 ));
  th24comp  U71_U_0_U_0 (.y ( f_n1_N_0 ) , .d ( f_n56 ) , .c ( t_n55 ) , .b ( f_n55 ) , .a ( t_n56 ));
  th24comp  U71_U_U (.y ( t_N7 ) , .d ( f_n1_N_0 ) , .c ( f_n54 ) , .b ( t_n54 ) , .a ( t_n1_N_0 ));
  th24comp  U71_U_U_0 (.y ( f_N7 ) , .d ( f_n1_N_0 ) , .c ( t_n54 ) , .b ( f_n54 ) , .a ( t_n1_N_0 ));
  th24comp  U86_U_0_U (.y ( t_n1_N ) , .d ( f_shift2_reg[0] ) , .c ( f_mul_reg[7] ) , .b ( t_mul_reg[7] ) , .a ( t_shift2_reg[0] ));
  th24comp  U86_U_0_U_0 (.y ( f_n1_N ) , .d ( f_shift2_reg[0] ) , .c ( t_mul_reg[7] ) , .b ( f_mul_reg[7] ) , .a ( t_shift2_reg[0] ));
  th24comp  U86_U_U (.y ( t_N16 ) , .d ( f_n1_N ) , .c ( f_n77 ) , .b ( t_n77 ) , .a ( t_n1_N ));
  th24comp  U86_U_U_0 (.y ( f_N16 ) , .d ( f_n1_N ) , .c ( t_n77 ) , .b ( f_n77 ) , .a ( t_n1_N ));
  drlatn  shift2_reg_reg_0__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N ) , .ackin ( acknet38 ) , .f_d ( f_q2_N ) , .t_d ( t_q2_N ) , .f_q ( f_shift2_reg[0] ) , .t_q ( t_shift2_reg[0] ));
  drlatr  shift2_reg_reg_0__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N ) , .ackin ( n2_N ) , .f_d ( f_q1_N ) , .t_d ( t_q1_N ) , .f_q ( f_q2_N ) , .t_q ( t_q2_N ));
  drlatn  shift2_reg_reg_0__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet0 ) , .ackin ( n1_N ) , .f_d ( f_constnet0 ) , .t_d ( t_constnet0 ) , .f_q ( f_q1_N ) , .t_q ( t_q1_N ));
  drlatn  mac_out_reg_0__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_0 ) , .ackin ( bufnet_2 ) , .f_d ( f_q2_N_0 ) , .t_d ( t_q2_N_0 ) , .f_q ( f_mac_out[0] ) , .t_q ( t_mac_out[0] ));
  drlatr  mac_out_reg_0__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_0 ) , .ackin ( n2_N_0 ) , .f_d ( f_q1_N_0 ) , .t_d ( t_q1_N_0 ) , .f_q ( f_q2_N_0 ) , .t_q ( t_q2_N_0 ));
  drlatn  mac_out_reg_0__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet1 ) , .ackin ( n1_N_0 ) , .f_d ( f_N9 ) , .t_d ( t_N9 ) , .f_q ( f_q1_N_0 ) , .t_q ( t_q1_N_0 ));
  drlatn  mac_out_reg_1__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_1 ) , .ackin ( bufnet_2 ) , .f_d ( f_q2_N_1 ) , .t_d ( t_q2_N_1 ) , .f_q ( f_mac_out[1] ) , .t_q ( t_mac_out[1] ));
  drlatr  mac_out_reg_1__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_1 ) , .ackin ( n2_N_1 ) , .f_d ( f_q1_N_1 ) , .t_d ( t_q1_N_1 ) , .f_q ( f_q2_N_1 ) , .t_q ( t_q2_N_1 ));
  drlatn  mac_out_reg_1__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet2 ) , .ackin ( n1_N_1 ) , .f_d ( f_N10 ) , .t_d ( t_N10 ) , .f_q ( f_q1_N_1 ) , .t_q ( t_q1_N_1 ));
  drlatn  mac_out_reg_2__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_2 ) , .ackin ( bufnet_2 ) , .f_d ( f_q2_N_2 ) , .t_d ( t_q2_N_2 ) , .f_q ( f_mac_out[2] ) , .t_q ( t_mac_out[2] ));
  drlatr  mac_out_reg_2__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_2 ) , .ackin ( n2_N_2 ) , .f_d ( f_q1_N_2 ) , .t_d ( t_q1_N_2 ) , .f_q ( f_q2_N_2 ) , .t_q ( t_q2_N_2 ));
  drlatn  mac_out_reg_2__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet3 ) , .ackin ( n1_N_2 ) , .f_d ( f_N11 ) , .t_d ( t_N11 ) , .f_q ( f_q1_N_2 ) , .t_q ( t_q1_N_2 ));
  drlatn  mac_out_reg_3__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_3 ) , .ackin ( bufnet_2 ) , .f_d ( f_q2_N_3 ) , .t_d ( t_q2_N_3 ) , .f_q ( f_mac_out[3] ) , .t_q ( t_mac_out[3] ));
  drlatr  mac_out_reg_3__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_3 ) , .ackin ( n2_N_3 ) , .f_d ( f_q1_N_3 ) , .t_d ( t_q1_N_3 ) , .f_q ( f_q2_N_3 ) , .t_q ( t_q2_N_3 ));
  drlatn  mac_out_reg_3__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet4 ) , .ackin ( n1_N_3 ) , .f_d ( f_N12 ) , .t_d ( t_N12 ) , .f_q ( f_q1_N_3 ) , .t_q ( t_q1_N_3 ));
  drlatn  mac_out_reg_4__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_4 ) , .ackin ( bufnet_2 ) , .f_d ( f_q2_N_4 ) , .t_d ( t_q2_N_4 ) , .f_q ( f_mac_out[4] ) , .t_q ( t_mac_out[4] ));
  drlatr  mac_out_reg_4__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_4 ) , .ackin ( n2_N_4 ) , .f_d ( f_q1_N_4 ) , .t_d ( t_q1_N_4 ) , .f_q ( f_q2_N_4 ) , .t_q ( t_q2_N_4 ));
  drlatn  mac_out_reg_4__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet5 ) , .ackin ( n1_N_4 ) , .f_d ( f_N13 ) , .t_d ( t_N13 ) , .f_q ( f_q1_N_4 ) , .t_q ( t_q1_N_4 ));
  drlatn  mac_out_reg_5__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_5 ) , .ackin ( bufnet_2 ) , .f_d ( f_q2_N_5 ) , .t_d ( t_q2_N_5 ) , .f_q ( f_mac_out[5] ) , .t_q ( t_mac_out[5] ));
  drlatr  mac_out_reg_5__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_5 ) , .ackin ( n2_N_5 ) , .f_d ( f_q1_N_5 ) , .t_d ( t_q1_N_5 ) , .f_q ( f_q2_N_5 ) , .t_q ( t_q2_N_5 ));
  drlatn  mac_out_reg_5__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet6 ) , .ackin ( n1_N_5 ) , .f_d ( f_N14 ) , .t_d ( t_N14 ) , .f_q ( f_q1_N_5 ) , .t_q ( t_q1_N_5 ));
  drlatn  mac_out_reg_6__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_6 ) , .ackin ( bufnet_2 ) , .f_d ( f_q2_N_6 ) , .t_d ( t_q2_N_6 ) , .f_q ( f_mac_out[6] ) , .t_q ( t_mac_out[6] ));
  drlatr  mac_out_reg_6__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_6 ) , .ackin ( n2_N_6 ) , .f_d ( f_q1_N_6 ) , .t_d ( t_q1_N_6 ) , .f_q ( f_q2_N_6 ) , .t_q ( t_q2_N_6 ));
  drlatn  mac_out_reg_6__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet7 ) , .ackin ( n1_N_6 ) , .f_d ( f_N15 ) , .t_d ( t_N15 ) , .f_q ( f_q1_N_6 ) , .t_q ( t_q1_N_6 ));
  drlatn  mac_out_reg_7__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_7 ) , .ackin ( bufnet_2 ) , .f_d ( f_q2_N_7 ) , .t_d ( t_q2_N_7 ) , .f_q ( f_mac_out[7] ) , .t_q ( t_mac_out[7] ));
  drlatr  mac_out_reg_7__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_7 ) , .ackin ( n2_N_7 ) , .f_d ( f_q1_N_7 ) , .t_d ( t_q1_N_7 ) , .f_q ( f_q2_N_7 ) , .t_q ( t_q2_N_7 ));
  drlatn  mac_out_reg_7__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet8 ) , .ackin ( n1_N_7 ) , .f_d ( f_N16 ) , .t_d ( t_N16 ) , .f_q ( f_q1_N_7 ) , .t_q ( t_q1_N_7 ));
  drlatn  shift2_reg_reg_1__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_8 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_8 ) , .t_d ( t_q2_N_8 ) , .f_q ( f_shift2_reg[1] ) , .t_q ( t_shift2_reg[1] ));
  drlatr  shift2_reg_reg_1__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_8 ) , .ackin ( n2_N_8 ) , .f_d ( f_q1_N_8 ) , .t_d ( t_q1_N_8 ) , .f_q ( f_q2_N_8 ) , .t_q ( t_q2_N_8 ));
  drlatn  shift2_reg_reg_1__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet9 ) , .ackin ( n1_N_8 ) , .f_d ( f_coef_reg[0] ) , .t_d ( t_coef_reg[0] ) , .f_q ( f_q1_N_8 ) , .t_q ( t_q1_N_8 ));
  drlatn  shift2_reg_reg_2__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_9 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_9 ) , .t_d ( t_q2_N_9 ) , .f_q ( f_shift2_reg[2] ) , .t_q ( t_shift2_reg[2] ));
  drlatr  shift2_reg_reg_2__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_9 ) , .ackin ( n2_N_9 ) , .f_d ( f_q1_N_9 ) , .t_d ( t_q1_N_9 ) , .f_q ( f_q2_N_9 ) , .t_q ( t_q2_N_9 ));
  drlatn  shift2_reg_reg_2__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet10 ) , .ackin ( n1_N_9 ) , .f_d ( f_coef_reg[1] ) , .t_d ( t_coef_reg[1] ) , .f_q ( f_q1_N_9 ) , .t_q ( t_q1_N_9 ));
  drlatn  shift2_reg_reg_3__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_10 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_10 ) , .t_d ( t_q2_N_10 ) , .f_q ( f_shift2_reg[3] ) , .t_q ( t_shift2_reg[3] ));
  drlatr  shift2_reg_reg_3__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_10 ) , .ackin ( n2_N_10 ) , .f_d ( f_q1_N_10 ) , .t_d ( t_q1_N_10 ) , .f_q ( f_q2_N_10 ) , .t_q ( t_q2_N_10 ));
  drlatn  shift2_reg_reg_3__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet11 ) , .ackin ( n1_N_10 ) , .f_d ( f_coef_reg[2] ) , .t_d ( t_coef_reg[2] ) , .f_q ( f_q1_N_10 ) , .t_q ( t_q1_N_10 ));
  drlatn  shift2_reg_reg_4__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_11 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_11 ) , .t_d ( t_q2_N_11 ) , .f_q ( f_shift2_reg[4] ) , .t_q ( t_shift2_reg[4] ));
  drlatr  shift2_reg_reg_4__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_11 ) , .ackin ( n2_N_11 ) , .f_d ( f_q1_N_11 ) , .t_d ( t_q1_N_11 ) , .f_q ( f_q2_N_11 ) , .t_q ( t_q2_N_11 ));
  drlatn  shift2_reg_reg_4__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet12 ) , .ackin ( n1_N_11 ) , .f_d ( f_coef_reg[3] ) , .t_d ( t_coef_reg[3] ) , .f_q ( f_q1_N_11 ) , .t_q ( t_q1_N_11 ));
  drlatn  mul_reg_reg_0__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_12 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_12 ) , .t_d ( t_q2_N_12 ) , .f_q ( f_mul_reg[0] ) , .t_q ( t_mul_reg[0] ));
  drlatr  mul_reg_reg_0__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_12 ) , .ackin ( n2_N_12 ) , .f_d ( f_q1_N_12 ) , .t_d ( t_q1_N_12 ) , .f_q ( f_q2_N_12 ) , .t_q ( t_q2_N_12 ));
  drlatn  mul_reg_reg_0__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet13 ) , .ackin ( n1_N_12 ) , .f_d ( f_N1 ) , .t_d ( t_N1 ) , .f_q ( f_q1_N_12 ) , .t_q ( t_q1_N_12 ));
  drlatn  mul_reg_reg_1__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_13 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_13 ) , .t_d ( t_q2_N_13 ) , .f_q ( f_mul_reg[1] ) , .t_q ( t_mul_reg[1] ));
  drlatr  mul_reg_reg_1__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_13 ) , .ackin ( n2_N_13 ) , .f_d ( f_q1_N_13 ) , .t_d ( t_q1_N_13 ) , .f_q ( f_q2_N_13 ) , .t_q ( t_q2_N_13 ));
  drlatn  mul_reg_reg_1__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet14 ) , .ackin ( n1_N_13 ) , .f_d ( f_N2 ) , .t_d ( t_N2 ) , .f_q ( f_q1_N_13 ) , .t_q ( t_q1_N_13 ));
  drlatn  mul_reg_reg_2__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_14 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_14 ) , .t_d ( t_q2_N_14 ) , .f_q ( f_mul_reg[2] ) , .t_q ( t_mul_reg[2] ));
  drlatr  mul_reg_reg_2__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_14 ) , .ackin ( n2_N_14 ) , .f_d ( f_q1_N_14 ) , .t_d ( t_q1_N_14 ) , .f_q ( f_q2_N_14 ) , .t_q ( t_q2_N_14 ));
  drlatn  mul_reg_reg_2__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet15 ) , .ackin ( n1_N_14 ) , .f_d ( f_N3 ) , .t_d ( t_N3 ) , .f_q ( f_q1_N_14 ) , .t_q ( t_q1_N_14 ));
  drlatn  mul_reg_reg_3__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_15 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_15 ) , .t_d ( t_q2_N_15 ) , .f_q ( f_mul_reg[3] ) , .t_q ( t_mul_reg[3] ));
  drlatr  mul_reg_reg_3__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_15 ) , .ackin ( n2_N_15 ) , .f_d ( f_q1_N_15 ) , .t_d ( t_q1_N_15 ) , .f_q ( f_q2_N_15 ) , .t_q ( t_q2_N_15 ));
  drlatn  mul_reg_reg_3__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet16 ) , .ackin ( n1_N_15 ) , .f_d ( f_N4 ) , .t_d ( t_N4 ) , .f_q ( f_q1_N_15 ) , .t_q ( t_q1_N_15 ));
  drlatn  mul_reg_reg_4__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_16 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_16 ) , .t_d ( t_q2_N_16 ) , .f_q ( f_mul_reg[4] ) , .t_q ( t_mul_reg[4] ));
  drlatr  mul_reg_reg_4__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_16 ) , .ackin ( n2_N_16 ) , .f_d ( f_q1_N_16 ) , .t_d ( t_q1_N_16 ) , .f_q ( f_q2_N_16 ) , .t_q ( t_q2_N_16 ));
  drlatn  mul_reg_reg_4__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet17 ) , .ackin ( n1_N_16 ) , .f_d ( f_N5 ) , .t_d ( t_N5 ) , .f_q ( f_q1_N_16 ) , .t_q ( t_q1_N_16 ));
  drlatn  mul_reg_reg_5__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_17 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_17 ) , .t_d ( t_q2_N_17 ) , .f_q ( f_mul_reg[5] ) , .t_q ( t_mul_reg[5] ));
  drlatr  mul_reg_reg_5__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_17 ) , .ackin ( n2_N_17 ) , .f_d ( f_q1_N_17 ) , .t_d ( t_q1_N_17 ) , .f_q ( f_q2_N_17 ) , .t_q ( t_q2_N_17 ));
  drlatn  mul_reg_reg_5__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet18 ) , .ackin ( n1_N_17 ) , .f_d ( f_N6 ) , .t_d ( t_N6 ) , .f_q ( f_q1_N_17 ) , .t_q ( t_q1_N_17 ));
  drlatn  mul_reg_reg_6__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_18 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_18 ) , .t_d ( t_q2_N_18 ) , .f_q ( f_mul_reg[6] ) , .t_q ( t_mul_reg[6] ));
  drlatr  mul_reg_reg_6__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_18 ) , .ackin ( n2_N_18 ) , .f_d ( f_q1_N_18 ) , .t_d ( t_q1_N_18 ) , .f_q ( f_q2_N_18 ) , .t_q ( t_q2_N_18 ));
  drlatn  mul_reg_reg_6__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet19 ) , .ackin ( n1_N_18 ) , .f_d ( f_N7 ) , .t_d ( t_N7 ) , .f_q ( f_q1_N_18 ) , .t_q ( t_q1_N_18 ));
  drlatn  mul_reg_reg_7__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_19 ) , .ackin ( acknet38 ) , .f_d ( f_q2_N_19 ) , .t_d ( t_q2_N_19 ) , .f_q ( f_mul_reg[7] ) , .t_q ( t_mul_reg[7] ));
  drlatr  mul_reg_reg_7__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_19 ) , .ackin ( n2_N_19 ) , .f_d ( f_q1_N_19 ) , .t_d ( t_q1_N_19 ) , .f_q ( f_q2_N_19 ) , .t_q ( t_q2_N_19 ));
  drlatn  mul_reg_reg_7__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet20 ) , .ackin ( n1_N_19 ) , .f_d ( f_N8 ) , .t_d ( t_N8 ) , .f_q ( f_q1_N_19 ) , .t_q ( t_q1_N_19 ));
  drlatn  inb_reg_reg_0__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_20 ) , .ackin ( acknet35 ) , .f_d ( f_q2_N_20 ) , .t_d ( t_q2_N_20 ) , .f_q ( f_inb_reg[0] ) , .t_q ( t_inb_reg[0] ));
  drlatr  inb_reg_reg_0__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_20 ) , .ackin ( n2_N_20 ) , .f_d ( f_q1_N_20 ) , .t_d ( t_q1_N_20 ) , .f_q ( f_q2_N_20 ) , .t_q ( t_q2_N_20 ));
  drlatn  inb_reg_reg_0__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet21 ) , .ackin ( n1_N_20 ) , .f_d ( f_inb[0] ) , .t_d ( t_inb[0] ) , .f_q ( f_q1_N_20 ) , .t_q ( t_q1_N_20 ));
  drlatn  inb_reg_reg_1__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_21 ) , .ackin ( acknet35 ) , .f_d ( f_q2_N_21 ) , .t_d ( t_q2_N_21 ) , .f_q ( f_inb_reg[1] ) , .t_q ( t_inb_reg[1] ));
  drlatr  inb_reg_reg_1__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_21 ) , .ackin ( n2_N_21 ) , .f_d ( f_q1_N_21 ) , .t_d ( t_q1_N_21 ) , .f_q ( f_q2_N_21 ) , .t_q ( t_q2_N_21 ));
  drlatn  inb_reg_reg_1__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet22 ) , .ackin ( n1_N_21 ) , .f_d ( f_inb[1] ) , .t_d ( t_inb[1] ) , .f_q ( f_q1_N_21 ) , .t_q ( t_q1_N_21 ));
  drlatn  inb_reg_reg_2__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_22 ) , .ackin ( acknet35 ) , .f_d ( f_q2_N_22 ) , .t_d ( t_q2_N_22 ) , .f_q ( f_inb_reg[2] ) , .t_q ( t_inb_reg[2] ));
  drlatr  inb_reg_reg_2__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_22 ) , .ackin ( n2_N_22 ) , .f_d ( f_q1_N_22 ) , .t_d ( t_q1_N_22 ) , .f_q ( f_q2_N_22 ) , .t_q ( t_q2_N_22 ));
  drlatn  inb_reg_reg_2__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet23 ) , .ackin ( n1_N_22 ) , .f_d ( f_inb[2] ) , .t_d ( t_inb[2] ) , .f_q ( f_q1_N_22 ) , .t_q ( t_q1_N_22 ));
  drlatn  inb_reg_reg_3__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_23 ) , .ackin ( acknet35 ) , .f_d ( f_q2_N_23 ) , .t_d ( t_q2_N_23 ) , .f_q ( f_inb_reg[3] ) , .t_q ( t_inb_reg[3] ));
  drlatr  inb_reg_reg_3__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_23 ) , .ackin ( n2_N_23 ) , .f_d ( f_q1_N_23 ) , .t_d ( t_q1_N_23 ) , .f_q ( f_q2_N_23 ) , .t_q ( t_q2_N_23 ));
  drlatn  inb_reg_reg_3__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet24 ) , .ackin ( n1_N_23 ) , .f_d ( f_inb[3] ) , .t_d ( t_inb[3] ) , .f_q ( f_q1_N_23 ) , .t_q ( t_q1_N_23 ));
  drlatn  ina_reg_reg_0__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_24 ) , .ackin ( acknet35 ) , .f_d ( f_q2_N_24 ) , .t_d ( t_q2_N_24 ) , .f_q ( f_ina_reg[0] ) , .t_q ( t_ina_reg[0] ));
  drlatr  ina_reg_reg_0__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_24 ) , .ackin ( n2_N_24 ) , .f_d ( f_q1_N_24 ) , .t_d ( t_q1_N_24 ) , .f_q ( f_q2_N_24 ) , .t_q ( t_q2_N_24 ));
  drlatn  ina_reg_reg_0__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet25 ) , .ackin ( n1_N_24 ) , .f_d ( f_ina[0] ) , .t_d ( t_ina[0] ) , .f_q ( f_q1_N_24 ) , .t_q ( t_q1_N_24 ));
  drlatn  ina_reg_reg_1__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_25 ) , .ackin ( acknet35 ) , .f_d ( f_q2_N_25 ) , .t_d ( t_q2_N_25 ) , .f_q ( f_ina_reg[1] ) , .t_q ( t_ina_reg[1] ));
  drlatr  ina_reg_reg_1__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_25 ) , .ackin ( n2_N_25 ) , .f_d ( f_q1_N_25 ) , .t_d ( t_q1_N_25 ) , .f_q ( f_q2_N_25 ) , .t_q ( t_q2_N_25 ));
  drlatn  ina_reg_reg_1__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet26 ) , .ackin ( n1_N_25 ) , .f_d ( f_ina[1] ) , .t_d ( t_ina[1] ) , .f_q ( f_q1_N_25 ) , .t_q ( t_q1_N_25 ));
  drlatn  ina_reg_reg_2__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_26 ) , .ackin ( acknet35 ) , .f_d ( f_q2_N_26 ) , .t_d ( t_q2_N_26 ) , .f_q ( f_ina_reg[2] ) , .t_q ( t_ina_reg[2] ));
  drlatr  ina_reg_reg_2__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_26 ) , .ackin ( n2_N_26 ) , .f_d ( f_q1_N_26 ) , .t_d ( t_q1_N_26 ) , .f_q ( f_q2_N_26 ) , .t_q ( t_q2_N_26 ));
  drlatn  ina_reg_reg_2__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet27 ) , .ackin ( n1_N_26 ) , .f_d ( f_ina[2] ) , .t_d ( t_ina[2] ) , .f_q ( f_q1_N_26 ) , .t_q ( t_q1_N_26 ));
  drlatn  ina_reg_reg_3__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_27 ) , .ackin ( acknet35 ) , .f_d ( f_q2_N_27 ) , .t_d ( t_q2_N_27 ) , .f_q ( f_ina_reg[3] ) , .t_q ( t_ina_reg[3] ));
  drlatr  ina_reg_reg_3__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_27 ) , .ackin ( n2_N_27 ) , .f_d ( f_q1_N_27 ) , .t_d ( t_q1_N_27 ) , .f_q ( f_q2_N_27 ) , .t_q ( t_q2_N_27 ));
  drlatn  ina_reg_reg_3__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet28 ) , .ackin ( n1_N_27 ) , .f_d ( f_ina[3] ) , .t_d ( t_ina[3] ) , .f_q ( f_q1_N_27 ) , .t_q ( t_q1_N_27 ));
  drlatn  coef_reg_reg_0__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_28 ) , .ackin ( acknet9 ) , .f_d ( f_q2_N_28 ) , .t_d ( t_q2_N_28 ) , .f_q ( f_coef_reg[0] ) , .t_q ( t_coef_reg[0] ));
  drlatr  coef_reg_reg_0__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_28 ) , .ackin ( n2_N_28 ) , .f_d ( f_q1_N_28 ) , .t_d ( t_q1_N_28 ) , .f_q ( f_q2_N_28 ) , .t_q ( t_q2_N_28 ));
  drlatn  coef_reg_reg_0__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet29 ) , .ackin ( n1_N_28 ) , .f_d ( f_coef[0] ) , .t_d ( t_coef[0] ) , .f_q ( f_q1_N_28 ) , .t_q ( t_q1_N_28 ));
  drlatn  coef_reg_reg_1__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_29 ) , .ackin ( acknet10 ) , .f_d ( f_q2_N_29 ) , .t_d ( t_q2_N_29 ) , .f_q ( f_coef_reg[1] ) , .t_q ( t_coef_reg[1] ));
  drlatr  coef_reg_reg_1__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_29 ) , .ackin ( n2_N_29 ) , .f_d ( f_q1_N_29 ) , .t_d ( t_q1_N_29 ) , .f_q ( f_q2_N_29 ) , .t_q ( t_q2_N_29 ));
  drlatn  coef_reg_reg_1__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet30 ) , .ackin ( n1_N_29 ) , .f_d ( f_coef[1] ) , .t_d ( t_coef[1] ) , .f_q ( f_q1_N_29 ) , .t_q ( t_q1_N_29 ));
  drlatn  coef_reg_reg_2__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_30 ) , .ackin ( acknet11 ) , .f_d ( f_q2_N_30 ) , .t_d ( t_q2_N_30 ) , .f_q ( f_coef_reg[2] ) , .t_q ( t_coef_reg[2] ));
  drlatr  coef_reg_reg_2__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_30 ) , .ackin ( n2_N_30 ) , .f_d ( f_q1_N_30 ) , .t_d ( t_q1_N_30 ) , .f_q ( f_q2_N_30 ) , .t_q ( t_q2_N_30 ));
  drlatn  coef_reg_reg_2__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet31 ) , .ackin ( n1_N_30 ) , .f_d ( f_coef[2] ) , .t_d ( t_coef[2] ) , .f_q ( f_q1_N_30 ) , .t_q ( t_q1_N_30 ));
  drlatn  coef_reg_reg_3__0_U (.rsb ( bufnet_0 ) , .ackout ( n2_N_31 ) , .ackin ( acknet12 ) , .f_d ( f_q2_N_31 ) , .t_d ( t_q2_N_31 ) , .f_q ( f_coef_reg[3] ) , .t_q ( t_coef_reg[3] ));
  drlatr  coef_reg_reg_3__0_U_0 (.rsb ( bufnet_0 ) , .ackout ( n1_N_31 ) , .ackin ( n2_N_31 ) , .f_d ( f_q1_N_31 ) , .t_d ( t_q1_N_31 ) , .f_q ( f_q2_N_31 ) , .t_q ( t_q2_N_31 ));
  drlatn  coef_reg_reg_3__0_U_1 (.rsb ( bufnet_0 ) , .ackout ( acknet32 ) , .ackin ( n1_N_31 ) , .f_d ( f_coef[3] ) , .t_d ( t_coef[3] ) , .f_q ( f_q1_N_31 ) , .t_q ( t_q1_N_31 ));
  and2  constcell0_0_U (.y ( f_constnet0 ) , .b ( acknet0 ) , .a ( bufnet_0 ));
  logic_0  constcell0_0_U_0 (.y ( t_constnet0 ));
  inv4x  bufcomp (.a ( rst_n ) , .y ( bufnet ));
  inv8x  bufcomp_0 (.a ( bufnet ) , .y ( bufnet_0 ));
  inv4x  bufcomp_1 (.a ( ackin ) , .y ( bufnet_1 ));
  inv  bufcomp_2 (.y ( bufnet_2 ) , .a ( bufnet_1 ));
endmodule
